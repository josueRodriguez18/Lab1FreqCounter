//test bench for frequency counter
module test()